`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    Xor32bit 
//////////////////////////////////////////////////////////////////////////////////
module Xor32bit(
    input A,B,
    output ALUop6
    );
	 always @(A,B)
	begin
	 out_ALUop6 <= A ^ B;
	end
endmodule
