`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    FullAdder1bit
//////////////////////////////////////////////////////////////////////////////////
module FullAdder1bit(
    input A,FB,ALUop1_cin,
    output sum,cout
    );
assign sum=A^FB^ALUop1_cin;
assign cout=A&FB|FB&ALUop1_cin|ALUop1_cin&A;

endmodule
