module SignExtend (X, Y);
    input X;
    output[31:0] Y;

    begin
      assign Y[0] = X;
      assign Y[1] = X;
      assign Y[2] = X;
      assign Y[3] = X;
      assign Y[4] = X;
      assign Y[5] = X;
      assign Y[6] = X;
      assign Y[7] = X;
      assign Y[8] = X;
      assign Y[9] = X;
      assign Y[10] = X;
      assign Y[11] = X;
      assign Y[12] = X;
      assign Y[13] = X;
      assign Y[14] = X;
      assign Y[15] = X;
      assign Y[16] = X;
      assign Y[17] = X;
      assign Y[18] = X;
      assign Y[19] = X;
      assign Y[20] = X;
      assign Y[21] = X;
      assign Y[22] = X;
      assign Y[23] = X;
      assign Y[24] = X;
      assign Y[25] = X;
      assign Y[26] = X;
      assign Y[27] = X;
      assign Y[28] = X;
      assign Y[29] = X;
      assign Y[30] = X;
      assign Y[31] = X;
    end

endmodule // SignExtend
