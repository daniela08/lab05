`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    Not32bit 
//////////////////////////////////////////////////////////////////////////////////
module Not32bit(
    input X,
    output Y
    );
	always @*
	begin
	 Y <= ~X;
	end
endmodule
