`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    Logic
//////////////////////////////////////////////////////////////////////////////////
module Logic(A, B, ALUop, LogicOut);
    input[31:0] A,B;
    input[3:0] ALUop;
    output[31:0] LogicOut;


endmodule
