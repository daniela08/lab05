module SignExtend (X, Y);
    input X;
    output[31:0] Y;

    begin
    Y[0] = X;
    Y[1] = X;
    Y[2] = X;
    Y[3] = X;
    Y[4] = X;
    Y[5] = X;
    Y[6] = X;
    Y[7] = X;
    Y[8] = X;
    Y[9] = X;
    Y[10] = X;
    Y[11] = X;
    Y[12] = X;
    Y[13] = X;
    Y[14] = X;
    Y[15] = X;
    Y[16] = X;
    Y[17] = X;
    Y[18] = X;
    Y[19] = X;
    Y[20] = X;
    Y[21] = X;
    Y[22] = X;
    Y[23] = X;
    Y[24] = X;
    Y[25] = X;
    Y[26] = X;
    Y[27] = X;
    Y[28] = X;
    Y[29] = X;
    Y[30] = X;
    Y[31] = X;
    end

endmodule // SignExtend
