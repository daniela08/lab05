`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    Not32bit
//////////////////////////////////////////////////////////////////////////////////
module Not32bit(
    input[31:0] X,
    output reg[31:0] Y);
	always @*
	begin
	 Y <= ~X;
	end

endmodule
